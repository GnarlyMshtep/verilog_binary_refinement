


module tester(); //or test bench 

//registers )

endmodule